`default_nettype none

module skullfet_inverter(input wire A, output reg Y);
    assign Y = !A;
endmodule
