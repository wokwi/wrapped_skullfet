`default_nettype none

module skullfet_inverter(input wire A, output wire Y);
    assign Y = !A;
endmodule
