VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO skullfet_inverter
  CLASS BLOCK ;
  FOREIGN skullfet_inverter ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.500 BY 13.300 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT 0.550 8.150 5.750 13.300 ;
      LAYER li1 ;
        RECT 0.800 12.450 1.600 13.200 ;
        RECT 0.600 11.950 1.800 12.450 ;
      LAYER mcon ;
        RECT 0.700 12.050 1.000 12.350 ;
      LAYER met1 ;
        RECT 0.000 11.950 1.100 12.450 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT 0.550 0.000 5.750 5.700 ;
      LAYER li1 ;
        RECT 0.900 1.050 1.800 1.550 ;
        RECT 0.850 0.350 1.550 1.050 ;
      LAYER mcon ;
        RECT 1.000 1.150 1.300 1.450 ;
      LAYER met1 ;
        RECT 0.000 1.050 1.400 1.550 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.700800 ;
    PORT
      LAYER li1 ;
        RECT 0.000 10.550 1.500 11.050 ;
        RECT 0.000 2.950 0.500 10.550 ;
        RECT 0.000 2.450 1.600 2.950 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER li1 ;
        RECT 6.000 3.950 6.500 9.350 ;
    END
  END A
  OBS
      LAYER met1 ;
        RECT 0.610 8.380 1.420 8.650 ;
        RECT 4.930 8.380 5.740 8.650 ;
        RECT 0.340 7.840 1.690 8.380 ;
        RECT 4.660 7.840 6.010 8.380 ;
        RECT 0.610 7.570 2.230 7.840 ;
        RECT 4.120 7.570 5.740 7.840 ;
        RECT 1.420 7.300 2.500 7.570 ;
        RECT 3.850 7.300 4.930 7.570 ;
        RECT 1.960 7.030 3.040 7.300 ;
        RECT 3.310 7.030 4.390 7.300 ;
        RECT 2.500 6.490 3.850 7.030 ;
        RECT 1.960 6.220 3.040 6.490 ;
        RECT 3.310 6.220 4.390 6.490 ;
        RECT 0.610 5.950 2.500 6.220 ;
        RECT 3.850 5.950 6.010 6.220 ;
        RECT 0.340 5.680 1.960 5.950 ;
        RECT 4.390 5.680 6.010 5.950 ;
        RECT 0.340 5.410 1.420 5.680 ;
        RECT 4.930 5.410 6.010 5.680 ;
        RECT 0.340 5.140 1.150 5.410 ;
        RECT 5.200 5.140 6.010 5.410 ;
        RECT 0.610 4.870 0.880 5.140 ;
        RECT 5.470 4.870 5.740 5.140 ;
  END
END skullfet_inverter
END LIBRARY

