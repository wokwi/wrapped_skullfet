VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO skullfet_inverter
  CLASS BLOCK ;
  FOREIGN skullfet_inverter ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.700 BY 14.400 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT 3.050 8.750 8.250 13.900 ;
      LAYER li1 ;
        RECT 3.300 13.050 4.100 13.800 ;
        RECT 3.100 12.550 4.300 13.050 ;
      LAYER mcon ;
        RECT 3.200 12.650 3.500 12.950 ;
      LAYER met1 ;
        RECT 0.000 14.000 10.700 14.400 ;
        RECT 2.500 13.050 2.900 14.000 ;
        RECT 2.500 12.550 3.600 13.050 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT 3.050 0.600 8.250 6.300 ;
      LAYER li1 ;
        RECT 3.400 1.650 4.300 2.150 ;
        RECT 3.350 0.950 4.050 1.650 ;
      LAYER mcon ;
        RECT 3.500 1.750 3.800 2.050 ;
      LAYER met1 ;
        RECT 2.500 1.650 3.900 2.150 ;
        RECT 2.500 0.400 3.000 1.650 ;
        RECT 0.000 0.000 10.700 0.400 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.700800 ;
    PORT
      LAYER li1 ;
        RECT 2.500 11.150 4.000 11.650 ;
        RECT 2.500 3.550 3.000 11.150 ;
        RECT 2.500 3.050 4.100 3.550 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER li1 ;
        RECT 8.500 4.550 9.000 9.950 ;
    END
  END A
  OBS
      LAYER met1 ;
        RECT 3.110 8.980 3.920 9.250 ;
        RECT 7.430 8.980 8.240 9.250 ;
        RECT 2.840 8.440 4.190 8.980 ;
        RECT 7.160 8.440 8.510 8.980 ;
        RECT 3.110 8.170 4.730 8.440 ;
        RECT 6.620 8.170 8.240 8.440 ;
        RECT 3.920 7.900 5.000 8.170 ;
        RECT 6.350 7.900 7.430 8.170 ;
        RECT 4.460 7.630 5.540 7.900 ;
        RECT 5.810 7.630 6.890 7.900 ;
        RECT 5.000 7.090 6.350 7.630 ;
        RECT 4.460 6.820 5.540 7.090 ;
        RECT 5.810 6.820 6.890 7.090 ;
        RECT 3.110 6.550 5.000 6.820 ;
        RECT 6.350 6.550 8.510 6.820 ;
        RECT 2.840 6.280 4.460 6.550 ;
        RECT 6.890 6.280 8.510 6.550 ;
        RECT 2.840 6.010 3.920 6.280 ;
        RECT 7.430 6.010 8.510 6.280 ;
        RECT 2.840 5.740 3.650 6.010 ;
        RECT 7.700 5.740 8.510 6.010 ;
        RECT 3.110 5.470 3.380 5.740 ;
        RECT 7.970 5.470 8.240 5.740 ;
  END
END skullfet_inverter
END LIBRARY

