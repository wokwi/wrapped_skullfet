(* blackbox *)
module skullfet_inverter(A, Y);
    input A;
    output Y;
endmodule
