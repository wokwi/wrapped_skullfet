VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO skullfet_inverter
  CLASS BLOCK ;
  FOREIGN skullfet_inverter ;
  ORIGIN -0.200 14.050 ;
  SIZE 6.500 BY 13.300 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT 0.750 -5.900 5.950 -0.750 ;
      LAYER li1 ;
        RECT 1.000 -1.600 1.800 -0.850 ;
        RECT 0.800 -2.100 2.000 -1.600 ;
      LAYER mcon ;
        RECT 0.900 -2.000 1.200 -1.700 ;
      LAYER met1 ;
        RECT 0.200 -2.100 1.300 -1.600 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT 0.750 -14.050 5.950 -8.350 ;
      LAYER li1 ;
        RECT 1.100 -13.000 2.000 -12.500 ;
        RECT 1.050 -13.700 1.750 -13.000 ;
      LAYER mcon ;
        RECT 1.200 -12.900 1.500 -12.600 ;
      LAYER met1 ;
        RECT 0.200 -13.000 1.600 -12.500 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.700800 ;
    PORT
      LAYER li1 ;
        RECT 0.200 -3.500 1.700 -3.000 ;
        RECT 0.200 -11.100 0.700 -3.500 ;
        RECT 0.200 -11.600 1.800 -11.100 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER li1 ;
        RECT 6.200 -10.100 6.700 -4.700 ;
    END
  END A
  OBS
      LAYER met1 ;
        RECT 0.810 -5.670 1.620 -5.400 ;
        RECT 5.130 -5.670 5.940 -5.400 ;
        RECT 0.540 -6.210 1.890 -5.670 ;
        RECT 4.860 -6.210 6.210 -5.670 ;
        RECT 0.810 -6.480 2.430 -6.210 ;
        RECT 4.320 -6.480 5.940 -6.210 ;
        RECT 1.620 -6.750 2.700 -6.480 ;
        RECT 4.050 -6.750 5.130 -6.480 ;
        RECT 2.160 -7.020 3.240 -6.750 ;
        RECT 3.510 -7.020 4.590 -6.750 ;
        RECT 2.700 -7.560 4.050 -7.020 ;
        RECT 2.160 -7.830 3.240 -7.560 ;
        RECT 3.510 -7.830 4.590 -7.560 ;
        RECT 0.810 -8.100 2.700 -7.830 ;
        RECT 4.050 -8.100 6.210 -7.830 ;
        RECT 0.540 -8.370 2.160 -8.100 ;
        RECT 4.590 -8.370 6.210 -8.100 ;
        RECT 0.540 -8.640 1.620 -8.370 ;
        RECT 5.130 -8.640 6.210 -8.370 ;
        RECT 0.540 -8.910 1.350 -8.640 ;
        RECT 5.400 -8.910 6.210 -8.640 ;
        RECT 0.810 -9.180 1.080 -8.910 ;
        RECT 5.670 -9.180 5.940 -8.910 ;
  END
END skullfet_inverter
END LIBRARY

