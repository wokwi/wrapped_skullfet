VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO skullfet_inverter
  CLASS BLOCK ;
  FOREIGN skullfet_inverter ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.700 BY 14.400 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT 3.050 8.750 8.250 13.900 ;
      LAYER li1 ;
        RECT 3.300 13.050 4.100 13.800 ;
        RECT 3.100 12.550 4.300 13.050 ;
      LAYER mcon ;
        RECT 3.200 12.700 3.450 12.950 ;
      LAYER met1 ;
        RECT 0.000 14.000 10.700 14.400 ;
        RECT 2.500 13.050 2.900 14.000 ;
        RECT 2.500 12.600 3.500 13.050 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT 3.050 0.600 8.250 6.300 ;
      LAYER li1 ;
        RECT 3.400 1.650 4.300 2.150 ;
        RECT 3.350 0.950 4.050 1.650 ;
      LAYER mcon ;
        RECT 3.450 1.750 3.700 1.950 ;
      LAYER met1 ;
        RECT 2.500 1.650 3.750 2.050 ;
        RECT 2.500 0.400 3.000 1.650 ;
        RECT 0.000 0.000 10.700 0.400 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.700800 ;
    PORT
      LAYER li1 ;
        RECT 2.500 11.150 4.000 11.650 ;
        RECT 2.500 3.550 3.000 11.150 ;
        RECT 2.500 3.050 4.100 3.550 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER li1 ;
        RECT 8.500 4.550 9.000 9.950 ;
    END
  END A
  OBS
      LAYER met1 ;
        RECT 4.730 13.300 6.890 13.570 ;
        RECT 4.460 13.030 6.890 13.300 ;
        RECT 3.920 12.490 7.430 13.030 ;
        RECT 3.650 11.410 7.700 12.490 ;
        RECT 3.650 11.140 4.460 11.410 ;
        RECT 3.650 10.870 4.190 11.140 ;
        RECT 3.920 10.600 4.190 10.870 ;
        RECT 5.270 10.600 6.080 11.410 ;
        RECT 6.890 11.140 7.700 11.410 ;
        RECT 7.160 10.870 7.700 11.140 ;
        RECT 7.160 10.600 7.430 10.870 ;
        RECT 3.920 10.330 4.460 10.600 ;
        RECT 5.000 10.330 6.350 10.600 ;
        RECT 6.890 10.330 7.430 10.600 ;
        RECT 3.920 10.060 5.540 10.330 ;
        RECT 5.810 10.060 7.160 10.330 ;
        RECT 4.460 9.790 5.270 10.060 ;
        RECT 6.080 9.790 7.160 10.060 ;
        RECT 4.730 9.250 6.620 9.790 ;
        RECT 3.110 8.980 3.920 9.250 ;
        RECT 4.730 8.980 5.000 9.250 ;
        RECT 5.270 8.980 5.540 9.250 ;
        RECT 5.810 8.980 6.080 9.250 ;
        RECT 6.350 8.980 6.620 9.250 ;
        RECT 7.430 8.980 8.240 9.250 ;
        RECT 2.840 8.440 4.190 8.980 ;
        RECT 7.160 8.440 8.510 8.980 ;
        RECT 3.110 8.170 4.730 8.440 ;
        RECT 6.620 8.170 8.240 8.440 ;
        RECT 3.920 7.900 5.000 8.170 ;
        RECT 6.350 7.900 7.430 8.170 ;
        RECT 4.460 7.630 5.540 7.900 ;
        RECT 5.810 7.630 6.890 7.900 ;
        RECT 5.000 7.090 6.350 7.630 ;
        RECT 4.460 6.820 5.540 7.090 ;
        RECT 5.810 6.820 6.890 7.090 ;
        RECT 3.110 6.550 5.000 6.820 ;
        RECT 6.350 6.550 8.510 6.820 ;
        RECT 2.840 6.280 4.460 6.550 ;
        RECT 6.890 6.280 8.510 6.550 ;
        RECT 2.840 6.010 3.920 6.280 ;
        RECT 7.430 6.010 8.510 6.280 ;
        RECT 2.840 5.740 3.650 6.010 ;
        RECT 7.700 5.740 8.510 6.010 ;
        RECT 3.110 5.470 3.380 5.740 ;
        RECT 4.730 5.470 5.000 5.740 ;
        RECT 5.270 5.470 5.540 5.740 ;
        RECT 5.810 5.470 6.080 5.740 ;
        RECT 6.350 5.470 6.620 5.740 ;
        RECT 7.970 5.470 8.240 5.740 ;
        RECT 4.730 4.930 6.620 5.470 ;
        RECT 4.460 4.660 5.270 4.930 ;
        RECT 6.080 4.660 7.160 4.930 ;
        RECT 3.920 4.390 5.540 4.660 ;
        RECT 5.810 4.390 7.160 4.660 ;
        RECT 3.920 4.120 4.460 4.390 ;
        RECT 5.000 4.120 6.350 4.390 ;
        RECT 6.890 4.120 7.430 4.390 ;
        RECT 3.920 3.850 4.190 4.120 ;
        RECT 3.650 3.580 4.190 3.850 ;
        RECT 3.650 3.310 4.460 3.580 ;
        RECT 5.270 3.310 6.080 4.120 ;
        RECT 7.160 3.850 7.430 4.120 ;
        RECT 7.160 3.580 7.700 3.850 ;
        RECT 6.890 3.310 7.700 3.580 ;
        RECT 3.650 2.230 7.700 3.310 ;
        RECT 3.920 1.690 7.430 2.230 ;
        RECT 4.460 1.420 6.890 1.690 ;
        RECT 4.730 1.150 6.890 1.420 ;
  END
END skullfet_inverter
END LIBRARY

