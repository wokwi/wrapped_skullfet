VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO skullfet_nand
  CLASS BLOCK ;
  FOREIGN skullfet_nand ;
  ORIGIN 4.320 13.770 ;
  SIZE 15.660 BY 12.690 ;
  OBS
      LAYER nwell ;
        RECT 6.210 -8.640 11.340 -4.860 ;
        RECT 1.080 -9.720 11.340 -8.640 ;
        RECT 1.080 -13.770 5.670 -9.720 ;
      LAYER li1 ;
        RECT -2.295 -2.160 2.025 -1.620 ;
        RECT -2.295 -5.535 -1.755 -2.160 ;
        RECT 7.020 -2.970 9.720 -2.430 ;
        RECT 4.995 -3.645 6.750 -3.105 ;
        RECT 6.210 -4.185 9.045 -3.645 ;
        RECT 8.505 -5.535 9.045 -4.185 ;
        RECT -3.780 -12.960 -3.240 -8.505 ;
        RECT 8.505 -10.935 9.045 -8.775 ;
        RECT 4.995 -11.475 9.045 -10.935 ;
        RECT -2.970 -12.150 -0.270 -11.610 ;
        RECT 9.990 -12.420 10.530 -8.505 ;
        RECT 4.725 -12.960 10.530 -12.420 ;
      LAYER mcon ;
        RECT -3.645 -12.960 -3.240 -12.420 ;
        RECT 7.020 -12.960 7.425 -12.420 ;
      LAYER met1 ;
        RECT 0.810 -5.670 1.620 -5.400 ;
        RECT 5.130 -5.670 5.940 -5.400 ;
        RECT 0.540 -6.210 1.890 -5.670 ;
        RECT 4.860 -6.210 6.210 -5.670 ;
        RECT 0.810 -6.480 2.430 -6.210 ;
        RECT 4.320 -6.480 5.940 -6.210 ;
        RECT 1.620 -6.750 2.700 -6.480 ;
        RECT 4.050 -6.750 5.130 -6.480 ;
        RECT 2.160 -7.020 3.240 -6.750 ;
        RECT 3.510 -7.020 4.590 -6.750 ;
        RECT 2.700 -7.560 4.050 -7.020 ;
        RECT 2.160 -7.830 3.240 -7.560 ;
        RECT 3.510 -7.830 4.590 -7.560 ;
        RECT 0.810 -8.100 2.700 -7.830 ;
        RECT 4.050 -8.100 6.210 -7.830 ;
        RECT 0.540 -8.370 2.160 -8.100 ;
        RECT 4.590 -8.370 6.210 -8.100 ;
        RECT 0.540 -8.640 1.620 -8.370 ;
        RECT 5.130 -8.640 6.210 -8.370 ;
        RECT 0.540 -8.910 1.350 -8.640 ;
        RECT 5.400 -8.910 6.210 -8.640 ;
        RECT 0.810 -9.180 1.080 -8.910 ;
        RECT 5.670 -9.180 5.940 -8.910 ;
        RECT -3.780 -13.095 -1.620 -12.285 ;
        RECT 6.885 -13.230 10.935 -11.880 ;
  END
END skullfet_nand
END LIBRARY

